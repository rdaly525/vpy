module Foo(
  input [10:0] i0,
  output [11:0] o0,
  inout [2:0]  io0,
  input i1,
  output o1,
  inout io1
);

endmodule
